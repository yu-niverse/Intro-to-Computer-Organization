//Subject:      CO project 2 - Shift_Left_Two_32
//--------------------------------------------------------------------------------
//Version:     1
//--------------------------------------------------------------------------------
//--------------------------------------------------------------------------------
//Writer:      109550182
//----------------------------------------------
//Date:        2022/04/25
//----------------------------------------------
//Description: 
//--------------------------------------------------------------------------------
`timescale 1ns/1ps
module Shift_Left_Two_32(data_i, data_o);

//I/O ports                    
input [32-1:0] data_i;
output [32-1:0] data_o;

//Internal signals
wire [32-1:0] data_o;

//shift left 2
assign data_o = {data_i[29:0], 2'b00};

endmodule
